typedef uvm_sequencer#(my_transaction) my_sequencer;
// 定义一个my_sequencer类型，它是uvm_sequencer的一个实例，专门用于处理my_transaction类型的事务。
