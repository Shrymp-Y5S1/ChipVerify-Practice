module PC_Reg (
    input clk,
    input rst_sync,
    input stall_n,   // 0: stall, 1: work
    input flush,

    input        [31:0] jump_addr,
    input               jump,
    output logic [31:0] pc          // PC address for instruction fetch
);

  always_ff @(posedge clk) begin
    if (rst_sync) begin
      pc <= 0;
    end else if (flush) begin
      pc <= 0;
    end else if (jump) begin
      pc <= jump_addr;
    end else if (stall_n) begin
      pc <= pc + 3'h4;
    end
  end

endmodule
