package axi_pkg;
    parameter ID_WIDTH   = 4;
    parameter ADDR_WIDTH = 32;
endpackage
