package axi_pkg;
    parameter ID_WIDTH   = 4;
    parameter ADDR_WIDTH = 32;
    parameter DATA_WIDTH = 64;

    parameter FIXED = 2'b0;
    parameter INCR  = 2'b1;
    parameter WRAP  = 2'b10;

endpackage
